
module booth_mult_8bit_DW01_add_0 ( A, B, CI, SUM, CO );
  input [15:0] A;
  input [15:0] B;
  output [15:0] SUM;
  input CI;
  output CO;
  wire   n1;
  wire   [15:1] carry;
  assign SUM[3] = B[3];
  assign SUM[2] = B[2];
  assign SUM[1] = B[1];
  assign SUM[0] = B[0];

  FAX1 U1_15 ( .A(A[15]), .B(B[15]), .C(carry[15]), .YS(SUM[15]) );
  FAX1 U1_14 ( .A(A[14]), .B(B[14]), .C(carry[14]), .YC(carry[15]), .YS(
        SUM[14]) );
  FAX1 U1_13 ( .A(A[13]), .B(B[13]), .C(carry[13]), .YC(carry[14]), .YS(
        SUM[13]) );
  FAX1 U1_12 ( .A(A[12]), .B(B[12]), .C(carry[12]), .YC(carry[13]), .YS(
        SUM[12]) );
  FAX1 U1_11 ( .A(A[11]), .B(B[11]), .C(carry[11]), .YC(carry[12]), .YS(
        SUM[11]) );
  FAX1 U1_10 ( .A(A[10]), .B(B[10]), .C(carry[10]), .YC(carry[11]), .YS(
        SUM[10]) );
  FAX1 U1_9 ( .A(A[9]), .B(B[9]), .C(carry[9]), .YC(carry[10]), .YS(SUM[9]) );
  FAX1 U1_8 ( .A(A[8]), .B(B[8]), .C(carry[8]), .YC(carry[9]), .YS(SUM[8]) );
  FAX1 U1_7 ( .A(A[7]), .B(B[7]), .C(carry[7]), .YC(carry[8]), .YS(SUM[7]) );
  FAX1 U1_6 ( .A(A[6]), .B(B[6]), .C(carry[6]), .YC(carry[7]), .YS(SUM[6]) );
  FAX1 U1_5 ( .A(A[5]), .B(B[5]), .C(n1), .YC(carry[6]), .YS(SUM[5]) );
  AND2X1 U1 ( .A(B[4]), .B(A[4]), .Y(n1) );
  XOR2X1 U2 ( .A(B[4]), .B(A[4]), .Y(SUM[4]) );
endmodule


module booth_mult_8bit ( a, b, prod );
  input [7:0] a;
  input [7:0] b;
  output [15:0] prod;
  wire   \pp[3][15] , \pp[3][14] , \pp[3][13] , \pp[3][12] , \pp[3][11] ,
         \pp[3][10] , \pp[3][9] , \pp[3][8] , \pp[3][7] , \pp[3][6] ,
         \pp[2][15] , \pp[2][12] , \pp[2][11] , \pp[2][10] , \pp[2][9] ,
         \pp[2][8] , \pp[2][7] , \pp[2][6] , \pp[1][15] , \pp[1][10] ,
         \pp[1][9] , \pp[1][8] , \pp[1][7] , \pp[1][6] , \pp[1][5] ,
         \pp[1][4] , \pp[1][3] , \pp[1][2] , \pp[0][9] , \pp[0][8] ,
         \pp[0][7] , \pp[0][6] , \pp[0][5] , \pp[0][4] , \pp[0][3] ,
         \pp[0][2] , N48, N49, N50, N51, N52, N53, N54, N55, N56, N58, N59,
         N60, N61, N62, N63, N64, N65, N91, N92, N93, N94, N95, N96, N97, N98,
         N102, N103, N104, N105, N106, N107, N108, N109, N137, N138, N139,
         N140, N141, N142, N143, N144, N150, N151, N152, N153, N154, N155,
         N156, N157, N188, N189, N190, N191, N192, N193, N194, N195, N203,
         N204, N205, N206, N207, N208, N209, N210, n59, n60, n61, n62, n68,
         n69, n70, n71, n72, n73, n75, n76, n77, n78, n82, n83, n84, n85, n86,
         n87, n89, n90, n91, n92, n94, n95, n96, n97, n98, n99, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, N242, N241, N240,
         N239, N238, N237, N236, N235, N234, N233, N232, N231, N226, N225,
         N224, N223, N222, N221, N220, N219, N218, N217, N216, N215, N214,
         N213, N212, N211, \sub_61/carry[14] , \sub_61/carry[13] ,
         \sub_61/carry[12] , \sub_61/carry[11] , \sub_61/carry[10] ,
         \sub_61/carry[9] , \sub_61/carry[8] , \sub_60/carry[15] ,
         \sub_60/carry[14] , \sub_60/carry[13] , \sub_60/carry[12] ,
         \sub_60/carry[11] , \sub_60/carry[10] , \sub_60/carry[9] ,
         \sub_52/carry[12] , \sub_52/carry[11] , \sub_52/carry[10] ,
         \sub_52/carry[9] , \sub_52/carry[8] , \sub_52/carry[7] ,
         \sub_52/carry[6] , \sub_51/carry[13] , \sub_51/carry[12] ,
         \sub_51/carry[11] , \sub_51/carry[10] , \sub_51/carry[9] ,
         \sub_51/carry[8] , \sub_51/carry[7] , \sub_43/carry[10] ,
         \sub_43/carry[9] , \sub_43/carry[8] , \sub_43/carry[7] ,
         \sub_43/carry[6] , \sub_43/carry[5] , \sub_43/carry[4] ,
         \sub_42/carry[11] , \sub_42/carry[10] , \sub_42/carry[9] ,
         \sub_42/carry[8] , \sub_42/carry[7] , \sub_42/carry[6] ,
         \sub_42/carry[5] , \sub_34/carry[8] , \sub_34/carry[7] ,
         \sub_34/carry[6] , \sub_34/carry[5] , \sub_34/carry[4] ,
         \sub_34/carry[3] , \sub_34/carry[2] , \sub_33/carry[9] ,
         \sub_33/carry[8] , \sub_33/carry[7] , \sub_33/carry[6] ,
         \sub_33/carry[5] , \sub_33/carry[4] , \sub_33/carry[3] ,
         \add_1_root_add_0_root_add_66_3/carry[15] ,
         \add_1_root_add_0_root_add_66_3/carry[14] ,
         \add_1_root_add_0_root_add_66_3/carry[13] ,
         \add_1_root_add_0_root_add_66_3/carry[12] ,
         \add_1_root_add_0_root_add_66_3/carry[11] ,
         \add_1_root_add_0_root_add_66_3/carry[10] ,
         \add_1_root_add_0_root_add_66_3/carry[9] ,
         \add_1_root_add_0_root_add_66_3/carry[8] ,
         \add_1_root_add_0_root_add_66_3/carry[7] ,
         \add_1_root_add_0_root_add_66_3/carry[6] ,
         \add_1_root_add_0_root_add_66_3/carry[5] ,
         \add_1_root_add_0_root_add_66_3/carry[4] ,
         \add_1_root_add_0_root_add_66_3/carry[3] ,
         \add_2_root_add_0_root_add_66_3/carry[15] ,
         \add_2_root_add_0_root_add_66_3/carry[14] ,
         \add_2_root_add_0_root_add_66_3/carry[13] ,
         \add_2_root_add_0_root_add_66_3/carry[12] ,
         \add_2_root_add_0_root_add_66_3/carry[11] ,
         \add_2_root_add_0_root_add_66_3/carry[10] ,
         \add_2_root_add_0_root_add_66_3/carry[9] ,
         \add_2_root_add_0_root_add_66_3/carry[8] ,
         \add_2_root_add_0_root_add_66_3/carry[7] , n182, n183, n184, n185,
         n186, n187, n188, n189, n190, n191, n192, n193, n194, n195, n196,
         n197, n198, n199, n200, n201, n202, n203, n204, n205, n206, n207,
         n208, n209, n210, n211, n212, n213, n214, n215, n216, n217, n218,
         n219, n220, n221, n222, n223, n224, n225, n226, n227, n228, n229,
         n230, n231, n232, n233, n234, n235, n236, n237, n238, n239, n240,
         n241, n242, n243, n244, n245, n246, n247, n248, n249, n250, n251,
         n252, n253, n254, n255, n256, n257, n258, n259, n260, n261, n262,
         n263, n264, n265, n266, n267, n268, n269, n270, n271, n272, n273,
         n274, n275, n276, n277, n278, n279, n280, n281, n282, n283, n284,
         n285, n286, n287, n288, n289, n290, n291, n292, n293, n294, n295,
         n296, n297, n298, n299, n300, n301, n302, n303, n304, n305, n306,
         n307, n308, n309, n310, n311, n312;
  assign N48 = a[0];

  OAI21X1 U41 ( .A(n222), .B(n302), .C(n215), .Y(\pp[3][6] ) );
  AOI21X1 U52 ( .A(n71), .B(a[7]), .C(n72), .Y(n68) );
  OAI21X1 U53 ( .A(n310), .B(b[7]), .C(n222), .Y(n71) );
  NOR3X1 U56 ( .A(b[5]), .B(b[6]), .C(n309), .Y(n62) );
  XOR2X1 U57 ( .A(b[6]), .B(b[5]), .Y(n73) );
  OAI21X1 U58 ( .A(n302), .B(n223), .C(n208), .Y(N231) );
  AOI21X1 U67 ( .A(n85), .B(a[7]), .C(n86), .Y(n82) );
  OAI21X1 U68 ( .A(n311), .B(b[5]), .C(n223), .Y(n85) );
  NOR3X1 U71 ( .A(b[3]), .B(b[4]), .C(n310), .Y(n78) );
  XOR2X1 U72 ( .A(b[4]), .B(b[3]), .Y(n87) );
  OAI21X1 U73 ( .A(n302), .B(n204), .C(n198), .Y(\pp[1][2] ) );
  AOI21X1 U80 ( .A(n97), .B(a[7]), .C(n98), .Y(n94) );
  OAI21X1 U81 ( .A(n312), .B(b[3]), .C(n204), .Y(n97) );
  NOR3X1 U84 ( .A(b[1]), .B(b[2]), .C(n311), .Y(n92) );
  XOR2X1 U85 ( .A(b[2]), .B(b[1]), .Y(n99) );
  OAI21X1 U88 ( .A(n301), .B(n225), .C(n209), .Y(\pp[0][7] ) );
  AOI22X1 U89 ( .A(N64), .B(n106), .C(N54), .D(n103), .Y(n105) );
  AOI22X1 U92 ( .A(N63), .B(n106), .C(N53), .D(n103), .Y(n107) );
  AOI22X1 U95 ( .A(N62), .B(n106), .C(N52), .D(n103), .Y(n109) );
  AOI22X1 U98 ( .A(N61), .B(n106), .C(N51), .D(n103), .Y(n111) );
  AOI22X1 U101 ( .A(N60), .B(n106), .C(N50), .D(n103), .Y(n113) );
  AOI22X1 U104 ( .A(N59), .B(n106), .C(N49), .D(n103), .Y(n115) );
  NAND2X1 U105 ( .A(n200), .B(n199), .Y(N212) );
  AOI22X1 U107 ( .A(N58), .B(n106), .C(N48), .D(n103), .Y(n117) );
  AOI21X1 U110 ( .A(a[7]), .B(n104), .C(n120), .Y(n101) );
  OAI21X1 U111 ( .A(n302), .B(n225), .C(n194), .Y(N211) );
  booth_mult_8bit_DW01_add_0 add_0_root_add_0_root_add_66_3 ( .A({N242, N241, 
        N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, 1'b0, 1'b0, 
        1'b0, 1'b0}), .B({N226, N225, N224, N223, N222, N221, N220, N219, N218, 
        N217, N216, N215, N214, N213, N212, N211}), .CI(1'b0), .SUM(prod) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_3  ( .A(\pp[1][3] ), .B(n224), .C(
        \add_1_root_add_0_root_add_66_3/carry[3] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[4] ), .YS(N214) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_4  ( .A(\pp[1][4] ), .B(n210), .C(
        \add_1_root_add_0_root_add_66_3/carry[4] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[5] ), .YS(N215) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_5  ( .A(\pp[1][5] ), .B(n205), .C(
        \add_1_root_add_0_root_add_66_3/carry[5] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[6] ), .YS(N216) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_6  ( .A(\pp[1][6] ), .B(n216), .C(
        \add_1_root_add_0_root_add_66_3/carry[6] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[7] ), .YS(N217) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_7  ( .A(\pp[1][7] ), .B(\pp[0][7] ), 
        .C(\add_1_root_add_0_root_add_66_3/carry[7] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[8] ), .YS(N218) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_8  ( .A(\pp[1][8] ), .B(n201), .C(
        \add_1_root_add_0_root_add_66_3/carry[8] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[9] ), .YS(N219) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_9  ( .A(\pp[1][9] ), .B(n226), .C(
        \add_1_root_add_0_root_add_66_3/carry[9] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[10] ), .YS(N220) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_10  ( .A(n211), .B(n226), .C(
        \add_1_root_add_0_root_add_66_3/carry[10] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[11] ), .YS(N221) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_11  ( .A(n220), .B(n226), .C(
        \add_1_root_add_0_root_add_66_3/carry[11] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[12] ), .YS(N222) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_12  ( .A(n220), .B(n226), .C(
        \add_1_root_add_0_root_add_66_3/carry[12] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[13] ), .YS(N223) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_13  ( .A(n220), .B(n226), .C(
        \add_1_root_add_0_root_add_66_3/carry[13] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[14] ), .YS(N224) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_14  ( .A(n220), .B(n226), .C(
        \add_1_root_add_0_root_add_66_3/carry[14] ), .YC(
        \add_1_root_add_0_root_add_66_3/carry[15] ), .YS(N225) );
  FAX1 \add_1_root_add_0_root_add_66_3/U1_15  ( .A(n220), .B(n226), .C(
        \add_1_root_add_0_root_add_66_3/carry[15] ), .YS(N226) );
  FAX1 \add_2_root_add_0_root_add_66_3/U1_7  ( .A(\pp[3][7] ), .B(\pp[2][7] ), 
        .C(\add_2_root_add_0_root_add_66_3/carry[7] ), .YC(
        \add_2_root_add_0_root_add_66_3/carry[8] ), .YS(N234) );
  FAX1 \add_2_root_add_0_root_add_66_3/U1_8  ( .A(\pp[3][8] ), .B(\pp[2][8] ), 
        .C(\add_2_root_add_0_root_add_66_3/carry[8] ), .YC(
        \add_2_root_add_0_root_add_66_3/carry[9] ), .YS(N235) );
  FAX1 \add_2_root_add_0_root_add_66_3/U1_9  ( .A(\pp[3][9] ), .B(\pp[2][9] ), 
        .C(\add_2_root_add_0_root_add_66_3/carry[9] ), .YC(
        \add_2_root_add_0_root_add_66_3/carry[10] ), .YS(N236) );
  FAX1 \add_2_root_add_0_root_add_66_3/U1_10  ( .A(\pp[3][10] ), .B(
        \pp[2][10] ), .C(\add_2_root_add_0_root_add_66_3/carry[10] ), .YC(
        \add_2_root_add_0_root_add_66_3/carry[11] ), .YS(N237) );
  FAX1 \add_2_root_add_0_root_add_66_3/U1_11  ( .A(\pp[3][11] ), .B(
        \pp[2][11] ), .C(\add_2_root_add_0_root_add_66_3/carry[11] ), .YC(
        \add_2_root_add_0_root_add_66_3/carry[12] ), .YS(N238) );
  FAX1 \add_2_root_add_0_root_add_66_3/U1_12  ( .A(\pp[3][12] ), .B(n191), .C(
        \add_2_root_add_0_root_add_66_3/carry[12] ), .YC(
        \add_2_root_add_0_root_add_66_3/carry[13] ), .YS(N239) );
  FAX1 \add_2_root_add_0_root_add_66_3/U1_13  ( .A(\pp[3][13] ), .B(n213), .C(
        \add_2_root_add_0_root_add_66_3/carry[13] ), .YC(
        \add_2_root_add_0_root_add_66_3/carry[14] ), .YS(N240) );
  FAX1 \add_2_root_add_0_root_add_66_3/U1_14  ( .A(n206), .B(n213), .C(
        \add_2_root_add_0_root_add_66_3/carry[14] ), .YC(
        \add_2_root_add_0_root_add_66_3/carry[15] ), .YS(N241) );
  FAX1 \add_2_root_add_0_root_add_66_3/U1_15  ( .A(n202), .B(n213), .C(
        \add_2_root_add_0_root_add_66_3/carry[15] ), .YS(N242) );
  AND2X1 U175 ( .A(n182), .B(n186), .Y(\pp[0][3] ) );
  AND2X1 U176 ( .A(n219), .B(n218), .Y(\pp[0][2] ) );
  AND2X1 U177 ( .A(n196), .B(n212), .Y(\pp[1][10] ) );
  AND2X1 U178 ( .A(n197), .B(n214), .Y(\pp[2][15] ) );
  AND2X1 U179 ( .A(n184), .B(n188), .Y(\pp[0][5] ) );
  AND2X1 U180 ( .A(n183), .B(n187), .Y(\pp[0][4] ) );
  AND2X1 U181 ( .A(n185), .B(n189), .Y(\pp[0][6] ) );
  AND2X1 U182 ( .A(n203), .B(n193), .Y(\pp[0][8] ) );
  AND2X1 U183 ( .A(n197), .B(n190), .Y(\pp[2][12] ) );
  AND2X1 U184 ( .A(n195), .B(n192), .Y(\pp[3][15] ) );
  AND2X1 U185 ( .A(n203), .B(n227), .Y(\pp[0][9] ) );
  AND2X1 U186 ( .A(n196), .B(n221), .Y(\pp[1][15] ) );
  AND2X1 U187 ( .A(n195), .B(n207), .Y(\pp[3][14] ) );
  AND2X1 U188 ( .A(n217), .B(\pp[1][2] ), .Y(
        \add_1_root_add_0_root_add_66_3/carry[3] ) );
  BUFX2 U189 ( .A(n113), .Y(n182) );
  BUFX2 U190 ( .A(n111), .Y(n183) );
  BUFX2 U191 ( .A(n109), .Y(n184) );
  BUFX2 U192 ( .A(n107), .Y(n185) );
  AND2X1 U193 ( .A(a[3]), .B(n104), .Y(n114) );
  INVX1 U194 ( .A(n114), .Y(n186) );
  AND2X1 U195 ( .A(a[4]), .B(n104), .Y(n112) );
  INVX1 U196 ( .A(n112), .Y(n187) );
  AND2X1 U197 ( .A(a[5]), .B(n104), .Y(n110) );
  INVX1 U198 ( .A(n110), .Y(n188) );
  AND2X1 U199 ( .A(a[6]), .B(n104), .Y(n108) );
  INVX1 U200 ( .A(n108), .Y(n189) );
  AND2X1 U201 ( .A(N143), .B(n78), .Y(n84) );
  INVX1 U202 ( .A(n84), .Y(n190) );
  INVX1 U203 ( .A(\pp[2][12] ), .Y(n191) );
  AND2X1 U204 ( .A(N195), .B(n62), .Y(n69) );
  INVX1 U205 ( .A(n69), .Y(n192) );
  AND2X1 U206 ( .A(N55), .B(n103), .Y(n102) );
  INVX1 U207 ( .A(n102), .Y(n193) );
  AND2X1 U208 ( .A(N48), .B(n106), .Y(n121) );
  INVX1 U209 ( .A(n121), .Y(n194) );
  BUFX2 U210 ( .A(n68), .Y(n195) );
  BUFX2 U211 ( .A(n94), .Y(n196) );
  BUFX2 U212 ( .A(n82), .Y(n197) );
  AND2X1 U213 ( .A(N48), .B(n91), .Y(n90) );
  INVX1 U214 ( .A(n90), .Y(n198) );
  AND2X1 U215 ( .A(a[1]), .B(n104), .Y(n118) );
  INVX1 U216 ( .A(n118), .Y(n199) );
  BUFX2 U217 ( .A(n117), .Y(n200) );
  INVX1 U218 ( .A(\pp[0][8] ), .Y(n201) );
  INVX1 U219 ( .A(\pp[3][15] ), .Y(n202) );
  BUFX2 U220 ( .A(n101), .Y(n203) );
  AND2X1 U221 ( .A(n99), .B(n311), .Y(n89) );
  INVX1 U222 ( .A(n89), .Y(n204) );
  INVX1 U223 ( .A(\pp[0][5] ), .Y(n205) );
  INVX1 U224 ( .A(\pp[3][14] ), .Y(n206) );
  AND2X1 U225 ( .A(N194), .B(n62), .Y(n70) );
  INVX1 U226 ( .A(n70), .Y(n207) );
  AND2X1 U227 ( .A(N48), .B(n77), .Y(n76) );
  INVX1 U228 ( .A(n76), .Y(n208) );
  BUFX2 U229 ( .A(n105), .Y(n209) );
  INVX1 U230 ( .A(\pp[0][4] ), .Y(n210) );
  INVX1 U231 ( .A(\pp[1][10] ), .Y(n211) );
  AND2X1 U232 ( .A(N97), .B(n92), .Y(n96) );
  INVX1 U233 ( .A(n96), .Y(n212) );
  INVX1 U234 ( .A(\pp[2][15] ), .Y(n213) );
  AND2X1 U235 ( .A(N144), .B(n78), .Y(n83) );
  INVX1 U236 ( .A(n83), .Y(n214) );
  AND2X1 U237 ( .A(N48), .B(n61), .Y(n60) );
  INVX1 U238 ( .A(n60), .Y(n215) );
  INVX1 U239 ( .A(\pp[0][6] ), .Y(n216) );
  INVX1 U240 ( .A(\pp[0][2] ), .Y(n217) );
  AND2X1 U241 ( .A(a[2]), .B(n104), .Y(n116) );
  INVX1 U242 ( .A(n116), .Y(n218) );
  BUFX2 U243 ( .A(n115), .Y(n219) );
  INVX1 U244 ( .A(\pp[1][15] ), .Y(n220) );
  AND2X1 U245 ( .A(N98), .B(n92), .Y(n95) );
  INVX1 U246 ( .A(n95), .Y(n221) );
  AND2X1 U247 ( .A(n73), .B(n309), .Y(n59) );
  INVX1 U248 ( .A(n59), .Y(n222) );
  AND2X1 U249 ( .A(n87), .B(n310), .Y(n75) );
  INVX1 U250 ( .A(n75), .Y(n223) );
  INVX1 U251 ( .A(\pp[0][3] ), .Y(n224) );
  AND2X1 U252 ( .A(b[0]), .B(n312), .Y(n104) );
  INVX1 U253 ( .A(n104), .Y(n225) );
  INVX1 U254 ( .A(\pp[0][9] ), .Y(n226) );
  AND2X1 U255 ( .A(N56), .B(n103), .Y(n119) );
  INVX1 U256 ( .A(n119), .Y(n227) );
  OR2X1 U257 ( .A(n255), .B(n259), .Y(n260) );
  XNOR2X1 U258 ( .A(n277), .B(b[3]), .Y(n228) );
  AND2X1 U259 ( .A(b[0]), .B(b[1]), .Y(n106) );
  OR2X1 U260 ( .A(n232), .B(n251), .Y(n252) );
  OR2X1 U261 ( .A(n278), .B(n297), .Y(n298) );
  OR2X1 U262 ( .A(n232), .B(n239), .Y(n240) );
  XNOR2X1 U263 ( .A(n300), .B(b[5]), .Y(n229) );
  XNOR2X1 U264 ( .A(n254), .B(b[1]), .Y(n230) );
  OR2X1 U265 ( .A(n232), .B(n236), .Y(n237) );
  OR2X1 U266 ( .A(n278), .B(n282), .Y(n283) );
  AND2X1 U267 ( .A(N109), .B(n91), .Y(n98) );
  AND2X1 U268 ( .A(N157), .B(n77), .Y(n86) );
  AND2X1 U269 ( .A(N210), .B(n61), .Y(n72) );
  AND2X1 U270 ( .A(N65), .B(n106), .Y(n120) );
  OR2X1 U271 ( .A(n312), .B(b[0]), .Y(n231) );
  INVX1 U272 ( .A(n231), .Y(n103) );
  OR2X1 U273 ( .A(n232), .B(n242), .Y(n243) );
  OR2X1 U274 ( .A(n232), .B(n245), .Y(n246) );
  OR2X1 U275 ( .A(n255), .B(n262), .Y(n263) );
  OR2X1 U276 ( .A(n278), .B(n279), .Y(n280) );
  OR2X1 U277 ( .A(n232), .B(n248), .Y(n249) );
  OR2X1 U278 ( .A(n255), .B(n265), .Y(n266) );
  OR2X1 U279 ( .A(n255), .B(n268), .Y(n269) );
  OR2X1 U280 ( .A(n278), .B(n285), .Y(n286) );
  OR2X1 U281 ( .A(n255), .B(n271), .Y(n272) );
  OR2X1 U282 ( .A(n278), .B(n288), .Y(n289) );
  OR2X1 U283 ( .A(n255), .B(n274), .Y(n275) );
  OR2X1 U284 ( .A(n278), .B(n291), .Y(n292) );
  OR2X1 U285 ( .A(n278), .B(n294), .Y(n295) );
  OR2X1 U286 ( .A(n232), .B(n233), .Y(n234) );
  OR2X1 U287 ( .A(n255), .B(n256), .Y(n257) );
  INVX1 U288 ( .A(a[7]), .Y(n301) );
  AND2X1 U289 ( .A(b[3]), .B(n99), .Y(n91) );
  AND2X1 U290 ( .A(b[5]), .B(n87), .Y(n77) );
  AND2X1 U291 ( .A(b[7]), .B(n73), .Y(n61) );
  INVX1 U292 ( .A(b[2]), .Y(n254) );
  INVX1 U293 ( .A(b[4]), .Y(n277) );
  INVX1 U294 ( .A(b[6]), .Y(n300) );
  INVX1 U295 ( .A(b[3]), .Y(n311) );
  INVX1 U296 ( .A(b[5]), .Y(n310) );
  INVX1 U297 ( .A(a[2]), .Y(n303) );
  INVX1 U298 ( .A(a[3]), .Y(n304) );
  INVX1 U299 ( .A(a[1]), .Y(n308) );
  INVX1 U300 ( .A(a[4]), .Y(n305) );
  INVX1 U301 ( .A(a[5]), .Y(n306) );
  INVX1 U302 ( .A(a[6]), .Y(n307) );
  INVX1 U303 ( .A(N48), .Y(n302) );
  INVX1 U304 ( .A(b[1]), .Y(n312) );
  INVX1 U305 ( .A(b[7]), .Y(n309) );
  XOR2X1 U306 ( .A(n254), .B(b[3]), .Y(n232) );
  MUX2X1 U307 ( .B(N48), .A(N48), .S(b[2]), .Y(n233) );
  MUX2X1 U308 ( .B(n234), .A(n235), .S(n230), .Y(\pp[1][3] ) );
  MUX2X1 U309 ( .B(N91), .A(a[1]), .S(b[2]), .Y(n236) );
  MUX2X1 U310 ( .B(n237), .A(n238), .S(n230), .Y(\pp[1][4] ) );
  MUX2X1 U311 ( .B(N92), .A(a[2]), .S(b[2]), .Y(n239) );
  MUX2X1 U312 ( .B(n240), .A(n241), .S(n230), .Y(\pp[1][5] ) );
  MUX2X1 U313 ( .B(N93), .A(a[3]), .S(b[2]), .Y(n242) );
  MUX2X1 U314 ( .B(n243), .A(n244), .S(n230), .Y(\pp[1][6] ) );
  MUX2X1 U315 ( .B(N94), .A(a[4]), .S(b[2]), .Y(n245) );
  MUX2X1 U316 ( .B(n246), .A(n247), .S(n230), .Y(\pp[1][7] ) );
  MUX2X1 U317 ( .B(N95), .A(a[5]), .S(b[2]), .Y(n248) );
  MUX2X1 U318 ( .B(n249), .A(n250), .S(n230), .Y(\pp[1][8] ) );
  MUX2X1 U319 ( .B(N96), .A(a[6]), .S(b[2]), .Y(n251) );
  MUX2X1 U320 ( .B(n252), .A(n253), .S(n230), .Y(\pp[1][9] ) );
  MUX2X1 U321 ( .B(a[1]), .A(N102), .S(b[3]), .Y(n235) );
  MUX2X1 U322 ( .B(a[2]), .A(N103), .S(b[3]), .Y(n238) );
  MUX2X1 U323 ( .B(a[3]), .A(N104), .S(b[3]), .Y(n241) );
  MUX2X1 U324 ( .B(a[4]), .A(N105), .S(b[3]), .Y(n244) );
  MUX2X1 U325 ( .B(a[5]), .A(N106), .S(b[3]), .Y(n247) );
  MUX2X1 U326 ( .B(a[6]), .A(N107), .S(b[3]), .Y(n250) );
  MUX2X1 U327 ( .B(a[7]), .A(N108), .S(b[3]), .Y(n253) );
  XOR2X1 U328 ( .A(n277), .B(b[5]), .Y(n255) );
  MUX2X1 U329 ( .B(N48), .A(N48), .S(b[4]), .Y(n256) );
  MUX2X1 U330 ( .B(n257), .A(n258), .S(n228), .Y(N232) );
  MUX2X1 U331 ( .B(N137), .A(a[1]), .S(b[4]), .Y(n259) );
  MUX2X1 U332 ( .B(n260), .A(n261), .S(n228), .Y(\pp[2][6] ) );
  MUX2X1 U333 ( .B(N138), .A(a[2]), .S(b[4]), .Y(n262) );
  MUX2X1 U334 ( .B(n263), .A(n264), .S(n228), .Y(\pp[2][7] ) );
  MUX2X1 U335 ( .B(N139), .A(a[3]), .S(b[4]), .Y(n265) );
  MUX2X1 U336 ( .B(n266), .A(n267), .S(n228), .Y(\pp[2][8] ) );
  MUX2X1 U337 ( .B(N140), .A(a[4]), .S(b[4]), .Y(n268) );
  MUX2X1 U338 ( .B(n269), .A(n270), .S(n228), .Y(\pp[2][9] ) );
  MUX2X1 U339 ( .B(N141), .A(a[5]), .S(b[4]), .Y(n271) );
  MUX2X1 U340 ( .B(n272), .A(n273), .S(n228), .Y(\pp[2][10] ) );
  MUX2X1 U341 ( .B(N142), .A(a[6]), .S(b[4]), .Y(n274) );
  MUX2X1 U342 ( .B(n275), .A(n276), .S(n228), .Y(\pp[2][11] ) );
  MUX2X1 U343 ( .B(a[1]), .A(N150), .S(b[5]), .Y(n258) );
  MUX2X1 U344 ( .B(a[2]), .A(N151), .S(b[5]), .Y(n261) );
  MUX2X1 U345 ( .B(a[3]), .A(N152), .S(b[5]), .Y(n264) );
  MUX2X1 U346 ( .B(a[4]), .A(N153), .S(b[5]), .Y(n267) );
  MUX2X1 U347 ( .B(a[5]), .A(N154), .S(b[5]), .Y(n270) );
  MUX2X1 U348 ( .B(a[6]), .A(N155), .S(b[5]), .Y(n273) );
  MUX2X1 U349 ( .B(a[7]), .A(N156), .S(b[5]), .Y(n276) );
  XOR2X1 U350 ( .A(n300), .B(b[7]), .Y(n278) );
  MUX2X1 U351 ( .B(N48), .A(N48), .S(b[6]), .Y(n279) );
  MUX2X1 U352 ( .B(n280), .A(n281), .S(n229), .Y(\pp[3][7] ) );
  MUX2X1 U353 ( .B(N188), .A(a[1]), .S(b[6]), .Y(n282) );
  MUX2X1 U354 ( .B(n283), .A(n284), .S(n229), .Y(\pp[3][8] ) );
  MUX2X1 U355 ( .B(N189), .A(a[2]), .S(b[6]), .Y(n285) );
  MUX2X1 U356 ( .B(n286), .A(n287), .S(n229), .Y(\pp[3][9] ) );
  MUX2X1 U357 ( .B(N190), .A(a[3]), .S(b[6]), .Y(n288) );
  MUX2X1 U358 ( .B(n289), .A(n290), .S(n229), .Y(\pp[3][10] ) );
  MUX2X1 U359 ( .B(N191), .A(a[4]), .S(b[6]), .Y(n291) );
  MUX2X1 U360 ( .B(n292), .A(n293), .S(n229), .Y(\pp[3][11] ) );
  MUX2X1 U361 ( .B(N192), .A(a[5]), .S(b[6]), .Y(n294) );
  MUX2X1 U362 ( .B(n295), .A(n296), .S(n229), .Y(\pp[3][12] ) );
  MUX2X1 U363 ( .B(N193), .A(a[6]), .S(b[6]), .Y(n297) );
  MUX2X1 U364 ( .B(n298), .A(n299), .S(n229), .Y(\pp[3][13] ) );
  MUX2X1 U365 ( .B(a[1]), .A(N203), .S(b[7]), .Y(n281) );
  MUX2X1 U366 ( .B(a[2]), .A(N204), .S(b[7]), .Y(n284) );
  MUX2X1 U367 ( .B(a[3]), .A(N205), .S(b[7]), .Y(n287) );
  MUX2X1 U368 ( .B(a[4]), .A(N206), .S(b[7]), .Y(n290) );
  MUX2X1 U369 ( .B(a[5]), .A(N207), .S(b[7]), .Y(n293) );
  MUX2X1 U370 ( .B(a[6]), .A(N208), .S(b[7]), .Y(n296) );
  MUX2X1 U371 ( .B(a[7]), .A(N209), .S(b[7]), .Y(n299) );
  XOR2X1 U372 ( .A(n217), .B(\pp[1][2] ), .Y(N213) );
  XOR2X1 U373 ( .A(n301), .B(\sub_33/carry[9] ), .Y(N56) );
  AND2X1 U374 ( .A(\sub_33/carry[8] ), .B(n301), .Y(\sub_33/carry[9] ) );
  XOR2X1 U375 ( .A(\sub_33/carry[8] ), .B(n301), .Y(N55) );
  AND2X1 U376 ( .A(\sub_33/carry[7] ), .B(n307), .Y(\sub_33/carry[8] ) );
  XOR2X1 U377 ( .A(\sub_33/carry[7] ), .B(n307), .Y(N54) );
  AND2X1 U378 ( .A(\sub_33/carry[6] ), .B(n306), .Y(\sub_33/carry[7] ) );
  XOR2X1 U379 ( .A(\sub_33/carry[6] ), .B(n306), .Y(N53) );
  AND2X1 U380 ( .A(\sub_33/carry[5] ), .B(n305), .Y(\sub_33/carry[6] ) );
  XOR2X1 U381 ( .A(\sub_33/carry[5] ), .B(n305), .Y(N52) );
  AND2X1 U382 ( .A(\sub_33/carry[4] ), .B(n304), .Y(\sub_33/carry[5] ) );
  XOR2X1 U383 ( .A(\sub_33/carry[4] ), .B(n304), .Y(N51) );
  AND2X1 U384 ( .A(\sub_33/carry[3] ), .B(n303), .Y(\sub_33/carry[4] ) );
  XOR2X1 U385 ( .A(\sub_33/carry[3] ), .B(n303), .Y(N50) );
  AND2X1 U386 ( .A(n302), .B(n308), .Y(\sub_33/carry[3] ) );
  XOR2X1 U387 ( .A(n302), .B(n308), .Y(N49) );
  XOR2X1 U388 ( .A(n301), .B(\sub_34/carry[8] ), .Y(N65) );
  AND2X1 U389 ( .A(\sub_34/carry[7] ), .B(n301), .Y(\sub_34/carry[8] ) );
  XOR2X1 U390 ( .A(\sub_34/carry[7] ), .B(n301), .Y(N64) );
  AND2X1 U391 ( .A(\sub_34/carry[6] ), .B(n307), .Y(\sub_34/carry[7] ) );
  XOR2X1 U392 ( .A(\sub_34/carry[6] ), .B(n307), .Y(N63) );
  AND2X1 U393 ( .A(\sub_34/carry[5] ), .B(n306), .Y(\sub_34/carry[6] ) );
  XOR2X1 U394 ( .A(\sub_34/carry[5] ), .B(n306), .Y(N62) );
  AND2X1 U395 ( .A(\sub_34/carry[4] ), .B(n305), .Y(\sub_34/carry[5] ) );
  XOR2X1 U396 ( .A(\sub_34/carry[4] ), .B(n305), .Y(N61) );
  AND2X1 U397 ( .A(\sub_34/carry[3] ), .B(n304), .Y(\sub_34/carry[4] ) );
  XOR2X1 U398 ( .A(\sub_34/carry[3] ), .B(n304), .Y(N60) );
  AND2X1 U399 ( .A(\sub_34/carry[2] ), .B(n303), .Y(\sub_34/carry[3] ) );
  XOR2X1 U400 ( .A(\sub_34/carry[2] ), .B(n303), .Y(N59) );
  AND2X1 U401 ( .A(n302), .B(n308), .Y(\sub_34/carry[2] ) );
  XOR2X1 U402 ( .A(n302), .B(n308), .Y(N58) );
  XOR2X1 U403 ( .A(n301), .B(\sub_42/carry[11] ), .Y(N98) );
  AND2X1 U404 ( .A(\sub_42/carry[10] ), .B(n301), .Y(\sub_42/carry[11] ) );
  XOR2X1 U405 ( .A(\sub_42/carry[10] ), .B(n301), .Y(N97) );
  AND2X1 U406 ( .A(\sub_42/carry[9] ), .B(n307), .Y(\sub_42/carry[10] ) );
  XOR2X1 U407 ( .A(\sub_42/carry[9] ), .B(n307), .Y(N96) );
  AND2X1 U408 ( .A(\sub_42/carry[8] ), .B(n306), .Y(\sub_42/carry[9] ) );
  XOR2X1 U409 ( .A(\sub_42/carry[8] ), .B(n306), .Y(N95) );
  AND2X1 U410 ( .A(\sub_42/carry[7] ), .B(n305), .Y(\sub_42/carry[8] ) );
  XOR2X1 U411 ( .A(\sub_42/carry[7] ), .B(n305), .Y(N94) );
  AND2X1 U412 ( .A(\sub_42/carry[6] ), .B(n304), .Y(\sub_42/carry[7] ) );
  XOR2X1 U413 ( .A(\sub_42/carry[6] ), .B(n304), .Y(N93) );
  AND2X1 U414 ( .A(\sub_42/carry[5] ), .B(n303), .Y(\sub_42/carry[6] ) );
  XOR2X1 U415 ( .A(\sub_42/carry[5] ), .B(n303), .Y(N92) );
  AND2X1 U416 ( .A(n302), .B(n308), .Y(\sub_42/carry[5] ) );
  XOR2X1 U417 ( .A(n302), .B(n308), .Y(N91) );
  XOR2X1 U418 ( .A(n301), .B(\sub_43/carry[10] ), .Y(N109) );
  AND2X1 U419 ( .A(\sub_43/carry[9] ), .B(n301), .Y(\sub_43/carry[10] ) );
  XOR2X1 U420 ( .A(\sub_43/carry[9] ), .B(n301), .Y(N108) );
  AND2X1 U421 ( .A(\sub_43/carry[8] ), .B(n307), .Y(\sub_43/carry[9] ) );
  XOR2X1 U422 ( .A(\sub_43/carry[8] ), .B(n307), .Y(N107) );
  AND2X1 U423 ( .A(\sub_43/carry[7] ), .B(n306), .Y(\sub_43/carry[8] ) );
  XOR2X1 U424 ( .A(\sub_43/carry[7] ), .B(n306), .Y(N106) );
  AND2X1 U425 ( .A(\sub_43/carry[6] ), .B(n305), .Y(\sub_43/carry[7] ) );
  XOR2X1 U426 ( .A(\sub_43/carry[6] ), .B(n305), .Y(N105) );
  AND2X1 U427 ( .A(\sub_43/carry[5] ), .B(n304), .Y(\sub_43/carry[6] ) );
  XOR2X1 U428 ( .A(\sub_43/carry[5] ), .B(n304), .Y(N104) );
  AND2X1 U429 ( .A(\sub_43/carry[4] ), .B(n303), .Y(\sub_43/carry[5] ) );
  XOR2X1 U430 ( .A(\sub_43/carry[4] ), .B(n303), .Y(N103) );
  AND2X1 U431 ( .A(n302), .B(n308), .Y(\sub_43/carry[4] ) );
  XOR2X1 U432 ( .A(n302), .B(n308), .Y(N102) );
  AND2X1 U433 ( .A(\pp[2][6] ), .B(\pp[3][6] ), .Y(
        \add_2_root_add_0_root_add_66_3/carry[7] ) );
  XOR2X1 U434 ( .A(\pp[2][6] ), .B(\pp[3][6] ), .Y(N233) );
  XOR2X1 U435 ( .A(n301), .B(\sub_51/carry[13] ), .Y(N144) );
  AND2X1 U436 ( .A(\sub_51/carry[12] ), .B(n301), .Y(\sub_51/carry[13] ) );
  XOR2X1 U437 ( .A(\sub_51/carry[12] ), .B(n301), .Y(N143) );
  AND2X1 U438 ( .A(\sub_51/carry[11] ), .B(n307), .Y(\sub_51/carry[12] ) );
  XOR2X1 U439 ( .A(\sub_51/carry[11] ), .B(n307), .Y(N142) );
  AND2X1 U440 ( .A(\sub_51/carry[10] ), .B(n306), .Y(\sub_51/carry[11] ) );
  XOR2X1 U441 ( .A(\sub_51/carry[10] ), .B(n306), .Y(N141) );
  AND2X1 U442 ( .A(\sub_51/carry[9] ), .B(n305), .Y(\sub_51/carry[10] ) );
  XOR2X1 U443 ( .A(\sub_51/carry[9] ), .B(n305), .Y(N140) );
  AND2X1 U444 ( .A(\sub_51/carry[8] ), .B(n304), .Y(\sub_51/carry[9] ) );
  XOR2X1 U445 ( .A(\sub_51/carry[8] ), .B(n304), .Y(N139) );
  AND2X1 U446 ( .A(\sub_51/carry[7] ), .B(n303), .Y(\sub_51/carry[8] ) );
  XOR2X1 U447 ( .A(\sub_51/carry[7] ), .B(n303), .Y(N138) );
  AND2X1 U448 ( .A(n302), .B(n308), .Y(\sub_51/carry[7] ) );
  XOR2X1 U449 ( .A(n302), .B(n308), .Y(N137) );
  XOR2X1 U450 ( .A(n301), .B(\sub_52/carry[12] ), .Y(N157) );
  AND2X1 U451 ( .A(\sub_52/carry[11] ), .B(n301), .Y(\sub_52/carry[12] ) );
  XOR2X1 U452 ( .A(\sub_52/carry[11] ), .B(n301), .Y(N156) );
  AND2X1 U453 ( .A(\sub_52/carry[10] ), .B(n307), .Y(\sub_52/carry[11] ) );
  XOR2X1 U454 ( .A(\sub_52/carry[10] ), .B(n307), .Y(N155) );
  AND2X1 U455 ( .A(\sub_52/carry[9] ), .B(n306), .Y(\sub_52/carry[10] ) );
  XOR2X1 U456 ( .A(\sub_52/carry[9] ), .B(n306), .Y(N154) );
  AND2X1 U457 ( .A(\sub_52/carry[8] ), .B(n305), .Y(\sub_52/carry[9] ) );
  XOR2X1 U458 ( .A(\sub_52/carry[8] ), .B(n305), .Y(N153) );
  AND2X1 U459 ( .A(\sub_52/carry[7] ), .B(n304), .Y(\sub_52/carry[8] ) );
  XOR2X1 U460 ( .A(\sub_52/carry[7] ), .B(n304), .Y(N152) );
  AND2X1 U461 ( .A(\sub_52/carry[6] ), .B(n303), .Y(\sub_52/carry[7] ) );
  XOR2X1 U462 ( .A(\sub_52/carry[6] ), .B(n303), .Y(N151) );
  AND2X1 U463 ( .A(n302), .B(n308), .Y(\sub_52/carry[6] ) );
  XOR2X1 U464 ( .A(n302), .B(n308), .Y(N150) );
  XOR2X1 U465 ( .A(n301), .B(\sub_60/carry[15] ), .Y(N195) );
  AND2X1 U466 ( .A(\sub_60/carry[14] ), .B(n301), .Y(\sub_60/carry[15] ) );
  XOR2X1 U467 ( .A(\sub_60/carry[14] ), .B(n301), .Y(N194) );
  AND2X1 U468 ( .A(\sub_60/carry[13] ), .B(n307), .Y(\sub_60/carry[14] ) );
  XOR2X1 U469 ( .A(\sub_60/carry[13] ), .B(n307), .Y(N193) );
  AND2X1 U470 ( .A(\sub_60/carry[12] ), .B(n306), .Y(\sub_60/carry[13] ) );
  XOR2X1 U471 ( .A(\sub_60/carry[12] ), .B(n306), .Y(N192) );
  AND2X1 U472 ( .A(\sub_60/carry[11] ), .B(n305), .Y(\sub_60/carry[12] ) );
  XOR2X1 U473 ( .A(\sub_60/carry[11] ), .B(n305), .Y(N191) );
  AND2X1 U474 ( .A(\sub_60/carry[10] ), .B(n304), .Y(\sub_60/carry[11] ) );
  XOR2X1 U475 ( .A(\sub_60/carry[10] ), .B(n304), .Y(N190) );
  AND2X1 U476 ( .A(\sub_60/carry[9] ), .B(n303), .Y(\sub_60/carry[10] ) );
  XOR2X1 U477 ( .A(\sub_60/carry[9] ), .B(n303), .Y(N189) );
  AND2X1 U478 ( .A(n302), .B(n308), .Y(\sub_60/carry[9] ) );
  XOR2X1 U479 ( .A(n302), .B(n308), .Y(N188) );
  XOR2X1 U480 ( .A(n301), .B(\sub_61/carry[14] ), .Y(N210) );
  AND2X1 U481 ( .A(\sub_61/carry[13] ), .B(n301), .Y(\sub_61/carry[14] ) );
  XOR2X1 U482 ( .A(\sub_61/carry[13] ), .B(n301), .Y(N209) );
  AND2X1 U483 ( .A(\sub_61/carry[12] ), .B(n307), .Y(\sub_61/carry[13] ) );
  XOR2X1 U484 ( .A(\sub_61/carry[12] ), .B(n307), .Y(N208) );
  AND2X1 U485 ( .A(\sub_61/carry[11] ), .B(n306), .Y(\sub_61/carry[12] ) );
  XOR2X1 U486 ( .A(\sub_61/carry[11] ), .B(n306), .Y(N207) );
  AND2X1 U487 ( .A(\sub_61/carry[10] ), .B(n305), .Y(\sub_61/carry[11] ) );
  XOR2X1 U488 ( .A(\sub_61/carry[10] ), .B(n305), .Y(N206) );
  AND2X1 U489 ( .A(\sub_61/carry[9] ), .B(n304), .Y(\sub_61/carry[10] ) );
  XOR2X1 U490 ( .A(\sub_61/carry[9] ), .B(n304), .Y(N205) );
  AND2X1 U491 ( .A(\sub_61/carry[8] ), .B(n303), .Y(\sub_61/carry[9] ) );
  XOR2X1 U492 ( .A(\sub_61/carry[8] ), .B(n303), .Y(N204) );
  AND2X1 U493 ( .A(n302), .B(n308), .Y(\sub_61/carry[8] ) );
  XOR2X1 U494 ( .A(n302), .B(n308), .Y(N203) );
endmodule

